module inst_mem
(
    input   [4:0]   A,
    output  [31:0]  RD
);

parameter MAX_INDEX = 32;

reg    [31:0]   im    [MAX_INDEX-1:0];

assign RD = im [A];

// Instruction example
initial begin
    im[0] = { 6'b001000, 5'd0, 5'd16, 16'd15  }; //addi $s0, $0, 15
    im[1] = { 6'b001000, 5'd0, 5'd17, 16'd25  }; //addi $s1, $0, 25
    im[2] = { 6'b001000, 5'd0, 5'd18, 16'd20  }; //addi $s2, $0, 20
    im[3] = { 6'b000000, 5'd16, 5'd17, 5'd8, 5'd0, 6'b100000  }; //add $t0, $s0, $s1 //40
    im[4] = { 6'b101011, 5'd0, 5'd8, 16'd0  }; //sw $t0, 0($0)
    im[5] = { 6'b000000, 5'd17, 5'd18, 5'd8, 5'd0, 6'b100010  }; //sub $t0, $s1, $s2 //5
    im[6] = { 6'b101011, 5'd0, 5'd8, 16'd1  }; //sw $t0, 1($0)
    im[7] = { 6'b000000, 5'd16, 5'd18, 5'd8, 5'd0, 6'b100010  }; //sub $t0, $s0, $s2 //-5
    im[8] = { 6'b101011, 5'd0, 5'd8, 16'd2  }; //sw $t0, 2($0)
    im[9] = { 6'b000000, 5'd16, 5'd17, 5'd8, 5'b00000, 6'b100100  }; //and $t0, $s0, $s1 //9
    im[10] = { 6'b101011, 5'd0, 5'd8, 16'd3  }; //sw $t0, 3($0)
    im[11] = { 6'b000000, 5'd17, 5'd18, 5'd8, 5'b00000, 6'b100101  }; //or $t0, $s1, $s2 //29
    im[12] = { 6'b101011, 5'd0, 5'd8, 16'd4  }; //sw $t0, 4($0)
    im[13] = { 6'b000000, 5'd17, 5'd18, 5'd8, 5'b00000, 6'b101010  }; //slt $t0, $s1, $s2 //0
    im[14] = { 6'b000000, 5'd18, 5'd17, 5'd8, 5'b00000, 6'b101010  }; //slt $t0, $s2, s1 //1
    im[15] = { 6'b000000, 5'd17, 5'd17, 5'd8, 5'b00000, 6'b101010  }; //slt $t0, $s1, $s1 //0
    im[16] = { 6'b100011, 5'd0, 5'd19, 16'd0  }; //lw $s3, 0($0)
    im[17] = { 6'b100011, 5'd0, 5'd20, 16'd1  }; //lw $s4, 1($0)
    im[18] = { 6'b100011, 5'd0, 5'd21, 16'd2  }; //lw $s5, 2($0)
    im[19] = { 6'b100011, 5'd0, 5'd22, 16'd3  }; //lw $s6, 3($0)
    im[20] = { 6'b100011, 5'd0, 5'd23, 16'd4  }; //lw $s7, 4($0)
end

endmodule
